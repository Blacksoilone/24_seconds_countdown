module alu (
    input alu_srca
    input alu_srcb
    
);
    
endmodule